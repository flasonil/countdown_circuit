// counter.sv